//
// sawp Wave ROM Table
//
module sawp_table(
  input [7:0] index,
  output [15:0] signal
);
parameter PERIOD = 256; // length of table

assign signal = sawp;
logic [15:0] sawp;
        
always_ff @(index)
begin
case(index)
	8'hff: sawp = 16'h3fff ;
	8'hfe: sawp = 16'h3fdf ;
	8'hfd: sawp = 16'h3ebf ;
	8'hfc: sawp = 16'h3e9f ;
	8'hfb: sawp = 16'h3d7f ;
	8'hfa: sawp = 16'h3d5f ;
	8'hf9: sawp = 16'h3c3f ;
	8'hf8: sawp = 16'h3c1f ;
	8'hf7: sawp = 16'h3bff ;
	8'hf6: sawp = 16'h3bdf ;
	8'hf5: sawp = 16'h3abf ;
	8'hf4: sawp = 16'h3a9f ;
	8'hf3: sawp = 16'h397f ;
	8'hf2: sawp = 16'h395f ;
	8'hf1: sawp = 16'h383f ;
	8'hf0: sawp = 16'h381f ;
	8'hef: sawp = 16'h37ff ;
	8'hee: sawp = 16'h37df ;
	8'hed: sawp = 16'h36bf ;
	8'hec: sawp = 16'h369f ;
	8'heb: sawp = 16'h357f ;
	8'hea: sawp = 16'h355f ;
	8'he9: sawp = 16'h343f ;
	8'he8: sawp = 16'h341f ;
	8'he7: sawp = 16'h33ff ;
	8'he6: sawp = 16'h33df ;
	8'he5: sawp = 16'h32bf ;
	8'he4: sawp = 16'h329f ;
	8'he3: sawp = 16'h317f ;
	8'he2: sawp = 16'h315f ;
	8'he1: sawp = 16'h303f ;
	8'he0: sawp = 16'h301f ;
	8'hdf: sawp = 16'h2fff ;
	8'hde: sawp = 16'h2fdf ;
	8'hdd: sawp = 16'h2ebf ;
	8'hdc: sawp = 16'h2e9f ;
	8'hdb: sawp = 16'h2d7f ;
	8'hda: sawp = 16'h2d5f ;
	8'hd9: sawp = 16'h2c3f ;
	8'hd8: sawp = 16'h2c1f ;
	8'hd7: sawp = 16'h2bff ;
	8'hd6: sawp = 16'h2bdf ;
	8'hd5: sawp = 16'h2abf ;
	8'hd4: sawp = 16'h2a9f ;
	8'hd3: sawp = 16'h297f ;
	8'hd2: sawp = 16'h295f ;
	8'hd1: sawp = 16'h283f ;
	8'hd0: sawp = 16'h281f ;
	8'hcf: sawp = 16'h27ff ;
	8'hce: sawp = 16'h27df ;
	8'hcd: sawp = 16'h26bf ;
	8'hcc: sawp = 16'h269f ;
	8'hcb: sawp = 16'h257f ;
	8'hca: sawp = 16'h255f ;
	8'hc9: sawp = 16'h243f ;
	8'hc8: sawp = 16'h241f ;
	8'hc7: sawp = 16'h23ff ;
	8'hc6: sawp = 16'h23df ;
	8'hc5: sawp = 16'h22bf ;
	8'hc4: sawp = 16'h229f ;
	8'hc3: sawp = 16'h217f ;
	8'hc2: sawp = 16'h215f ;
	8'hc1: sawp = 16'h203f ;
	8'hc0: sawp = 16'h201f ;
	8'hbf: sawp = 16'h1fff ;
	8'hbe: sawp = 16'h1fdf ;
	8'hbd: sawp = 16'h1ebf ;
	8'hbc: sawp = 16'h1e9f ;
	8'hbb: sawp = 16'h1d7f ;
	8'hba: sawp = 16'h1d5f ;
	8'hb9: sawp = 16'h1c3f ;
	8'hb8: sawp = 16'h1c1f ;
	8'hb7: sawp = 16'h1bff ;
	8'hb6: sawp = 16'h1bdf ;
	8'hb5: sawp = 16'h1abf ;
	8'hb4: sawp = 16'h1a9f ;
	8'hb3: sawp = 16'h197f ;
	8'hb2: sawp = 16'h195f ;
	8'hb1: sawp = 16'h183f ;
	8'hb0: sawp = 16'h181f ;
	8'haf: sawp = 16'h17ff ;
	8'hae: sawp = 16'h17df ;
	8'had: sawp = 16'h16bf ;
	8'hac: sawp = 16'h169f ;
	8'hab: sawp = 16'h157f ;
	8'haa: sawp = 16'h155f ;
	8'ha9: sawp = 16'h143f ;
	8'ha8: sawp = 16'h141f ;
	8'ha7: sawp = 16'h13ff ;
	8'ha6: sawp = 16'h13df ;
	8'ha5: sawp = 16'h12bf ;
	8'ha4: sawp = 16'h129f ;
	8'ha3: sawp = 16'h117f ;
	8'ha2: sawp = 16'h115f ;
	8'ha1: sawp = 16'h103f ;
	8'ha0: sawp = 16'h101f ;
	8'h9f: sawp = 16'h0fff ;
	8'h9e: sawp = 16'h0fdf ;
	8'h9d: sawp = 16'h0ebf ;
	8'h9c: sawp = 16'h0e9f ;
	8'h9b: sawp = 16'h0d7f ;
	8'h9a: sawp = 16'h0d5f ;
	8'h99: sawp = 16'h0c3f ;
	8'h98: sawp = 16'h0c1f ;
	8'h97: sawp = 16'h0bff ;
	8'h96: sawp = 16'h0bdf ;
	8'h95: sawp = 16'h0abf ;
	8'h94: sawp = 16'h0a9f ;
	8'h93: sawp = 16'h097f ;
	8'h92: sawp = 16'h095f ;
	8'h91: sawp = 16'h083f ;
	8'h90: sawp = 16'h081f ;
	8'h8f: sawp = 16'h07ff ;
	8'h8e: sawp = 16'h07df ;
	8'h8d: sawp = 16'h06bf ;
	8'h8c: sawp = 16'h069f ;
	8'h8b: sawp = 16'h057f ;
	8'h8a: sawp = 16'h0f5f ;
	8'h89: sawp = 16'h053f ;
	8'h88: sawp = 16'h041f ;
	8'h87: sawp = 16'h04ff ;
	8'h86: sawp = 16'h03df ;
	8'h85: sawp = 16'h03bf ;
	8'h84: sawp = 16'h029f ;
	8'h83: sawp = 16'h027f ;
	8'h82: sawp = 16'h015f ;
	8'h81: sawp = 16'h013f ;
	8'h80: sawp = 16'h001f ;
	8'h7f: sawp = 16'h0000 ;
	8'h7e: sawp = 16'hffe1 ;
	8'h7d: sawp = 16'hffc1 ;
	8'h7c: sawp = 16'hfea1 ;
	8'h7b: sawp = 16'hfe81 ;
	8'h7a: sawp = 16'hfd61 ;
	8'h79: sawp = 16'hfd41 ;
	8'h78: sawp = 16'hfc21 ;
	8'h77: sawp = 16'hfc01 ;
	8'h76: sawp = 16'hfbe1 ;
	8'h75: sawp = 16'hfbc1 ;
	8'h74: sawp = 16'hfaa1 ;
	8'h73: sawp = 16'hfa81 ;
	8'h72: sawp = 16'hf961 ;
	8'h71: sawp = 16'hf941 ;
	8'h70: sawp = 16'hf821 ;
	8'h6f: sawp = 16'hf801 ;
	8'h6e: sawp = 16'hf7e1 ;
	8'h6d: sawp = 16'hf7c1 ;
	8'h6c: sawp = 16'hf6a1 ;
	8'h6b: sawp = 16'hf681 ;
	8'h6a: sawp = 16'hf561 ;
	8'h69: sawp = 16'hf541 ;
	8'h68: sawp = 16'hf421 ;
	8'h67: sawp = 16'hf401 ;
	8'h66: sawp = 16'hf3e1 ;
	8'h65: sawp = 16'hf3c1 ;
	8'h64: sawp = 16'hf2a1 ;
	8'h63: sawp = 16'hf281 ;
	8'h62: sawp = 16'hf161 ;
	8'h61: sawp = 16'hf141 ;
	8'h60: sawp = 16'hf021 ;
	8'h5f: sawp = 16'hf001 ;
	8'h5e: sawp = 16'hefe1 ;
	8'h5d: sawp = 16'hefc1 ;
	8'h5c: sawp = 16'heea1 ;
	8'h5b: sawp = 16'hee81 ;
	8'h5a: sawp = 16'hed61 ;
	8'h59: sawp = 16'hed41 ;
	8'h58: sawp = 16'hec21 ;
	8'h57: sawp = 16'hec01 ;
	8'h56: sawp = 16'hebe1 ;
	8'h55: sawp = 16'hebc1 ;
	8'h54: sawp = 16'heaa1 ;
	8'h53: sawp = 16'hea81 ;
	8'h52: sawp = 16'he961 ;
	8'h51: sawp = 16'he941 ;
	8'h50: sawp = 16'he821 ;
	8'h4f: sawp = 16'he801 ;
	8'h4e: sawp = 16'he7e1 ;
	8'h4d: sawp = 16'he7c1 ;
	8'h4c: sawp = 16'he6a1 ;
	8'h4b: sawp = 16'he681 ;
	8'h4a: sawp = 16'he561 ;
	8'h49: sawp = 16'he541 ;
	8'h48: sawp = 16'he421 ;
	8'h47: sawp = 16'he401 ;
	8'h46: sawp = 16'he3e1 ;
	8'h45: sawp = 16'he3c1 ;
	8'h44: sawp = 16'he2a1 ;
	8'h43: sawp = 16'he281 ;
	8'h42: sawp = 16'he161 ;
	8'h41: sawp = 16'he141 ;
	8'h40: sawp = 16'he021 ;
	8'h3f: sawp = 16'he001 ;
	8'h3e: sawp = 16'hdfe1 ;
	8'h3d: sawp = 16'hdfc1 ;
	8'h3c: sawp = 16'hdea1 ;
	8'h3b: sawp = 16'hde81 ;
	8'h3a: sawp = 16'hdd61 ;
	8'h39: sawp = 16'hdd41 ;
	8'h38: sawp = 16'hdc21 ;
	8'h37: sawp = 16'hdc01 ;
	8'h36: sawp = 16'hdbe1 ;
	8'h35: sawp = 16'hdbc1 ;
	8'h34: sawp = 16'hdaa1 ;
	8'h33: sawp = 16'hda81 ;
	8'h32: sawp = 16'hd961 ;
	8'h31: sawp = 16'hd941 ;
	8'h30: sawp = 16'hd821 ;
	8'h2f: sawp = 16'hd801 ;
	8'h2e: sawp = 16'hd7e1 ;
	8'h2d: sawp = 16'hd7c1 ;
	8'h2c: sawp = 16'hd6a1 ;
	8'h2b: sawp = 16'hd681 ;
	8'h2a: sawp = 16'hd561 ;
	8'h29: sawp = 16'hd541 ;
	8'h28: sawp = 16'hd421 ;
	8'h27: sawp = 16'hd401 ;
	8'h26: sawp = 16'hd3e1 ;
	8'h25: sawp = 16'hd3c1 ;
	8'h24: sawp = 16'hd2a1 ;
	8'h23: sawp = 16'hd281 ;
	8'h22: sawp = 16'hd161 ;
	8'h21: sawp = 16'hd141 ;
	8'h20: sawp = 16'hd021 ;
	8'h1f: sawp = 16'hc001 ;
	8'h1e: sawp = 16'hcfe1 ;
	8'h1d: sawp = 16'hcfc1 ;
	8'h1c: sawp = 16'hcea1 ;
	8'h1b: sawp = 16'hce81 ;
	8'h1a: sawp = 16'hcd61 ;
	8'h19: sawp = 16'hcd41 ;
	8'h18: sawp = 16'hcc21 ;
	8'h17: sawp = 16'hcc01 ;
	8'h16: sawp = 16'hcbe1 ;
	8'h15: sawp = 16'hcbc1 ;
	8'h14: sawp = 16'hcaa1 ;
	8'h13: sawp = 16'hca81 ;
	8'h12: sawp = 16'hc961 ;
	8'h11: sawp = 16'hc941 ;
	8'h10: sawp = 16'hc821 ;
	8'h0f: sawp = 16'hc801 ;
	8'h0e: sawp = 16'hc7e1 ;
	8'h0d: sawp = 16'hc7c1 ;
	8'h0c: sawp = 16'hc6a1 ;
	8'h0b: sawp = 16'hc681 ;
	8'h0a: sawp = 16'hc561 ;
	8'h09: sawp = 16'hc541 ;
	8'h08: sawp = 16'hc421 ;
	8'h07: sawp = 16'hc401 ;
	8'h06: sawp = 16'hc3e1 ;
	8'h05: sawp = 16'hc3c1 ;
	8'h04: sawp = 16'hc2a1 ;
	8'h03: sawp = 16'hc281 ;
	8'h02: sawp = 16'hc161 ;
	8'h01: sawp = 16'hc141 ;
	8'h00: sawp = 16'hc021 ;
	default: sawp = 16'h0000;
endcase
end
endmodule
