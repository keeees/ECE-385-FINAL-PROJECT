module start(	input  frame_clk,Reset , 
					input [9:0] x,
					input [9:0] y,
					output logic [7:0] R,
					output logic [7:0] G,
					output logic [7:0] B
						);
	logic [2:0] pixel;
	logic [0:479][0:639][0:2] matrix;
	logic [5:0] counter;
	logic [2:0] cry;
	logic [2:0] tear,bkgd;
	
	 always_ff @ (posedge frame_clk)
    begin
        if (Reset)
        begin
            counter <= 6'd0;
				tear <= 3'd0;
				//cry <= 3'd0;
        end
        else
        begin
            counter <= counter +6'd1;
				if(counter <= 10'd12)
				tear <= 3'd2;
				//cry <= 3'd1;
				else if(counter > 6'd12 && counter <= 6'd24)
				tear <= 3'd3;
				//cry <= 3'd2;
				else if(counter > 6'd24 && counter <= 6'd36)
				tear <= 3'd4;
				//cry <= 3'd3;
				else if(counter > 6'd36 && counter <= 6'd48)
				tear <= 3'd5;
				//cry <= 3'd4;
				else if(counter > 6'd48 && counter <= 6'd60)
				tear <= 3'd6;
				//cry <= 3'd5;
				else counter <= 6'd0;
        end
    end


	
	always_comb begin
	

		  
		pixel = matrix[y-18][x];
		
		
		//tear = 3'd4;
		
		case(pixel)
		3'd0: begin
			R = 8'd255;
			G = 8'd255;
			B = 8'd255;

		end
		3'd1: begin//shen lv frog 
			R = 8'd0;
			G = 8'd95;
			B = 8'd29;
		end
		3'd2: begin//shen hong zuichun wai&press start
			R = 8'd149;
			G = 8'd23;
			B = 8'd0;
		end
		3'd3: begin//zuichun limian & xinyi gu
			R = 8'd255;
			G = 8'd129;
			B = 8'd117;
		end
		3'd4: begin// tears &sun ke
			R = 8'd60;
			G = 8'd241;
			B = 8'd255;
		end
		3'd5: begin //orange
			R = 8'd255;
			G = 8'd123;
			B = 8'd43;
		end
		3'd6: begin//yellow sun
			R = 8'd255;
			G = 8'd209;
			B = 8'd0;
		end
		3'd7: begin
			R = 8'd0;
			G = 8'd0;
			B = 8'd0;
		end
		bkgd:begin
		  R = 8'h3f; 
        G = 8'h00;
        B = 8'h7f - {1'b0, x[9:3]};
		end
		
		default:
		begin
		  R = 8'h3f; 
        G = 8'h00;
        B = 8'h7f - {1'b0, x[9:3]};
		  end
		  
		
		
		
	endcase
		
matrix = '{
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd5, 3'd5, 3'd5, 3'd5, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd4, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, tear, tear, tear, tear, tear, tear, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, tear, tear, tear, tear, tear, tear, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, tear, tear, tear, tear, tear, tear, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, tear, tear, tear, tear, tear, tear, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, tear, tear, tear, tear, tear, tear, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, tear, tear, tear, tear, tear, tear, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, tear, tear, tear, tear, tear, tear, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, tear, tear, tear, tear, tear, tear, tear, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, tear, tear, tear, tear, tear, tear, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd3, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, 3'd2, 3'd2, 3'd2, 3'd2, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd },
' {bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd, bkgd }

};
end
endmodule

















