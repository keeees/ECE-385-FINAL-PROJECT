module background(
					input [9:0] x,
					input [9:0] y,
					output logic [7:0] R,
					output logic [7:0] G,
					output logic [7:0] B
						);
	logic [1:0] pixel;
	logic [0:19][0:19][0:1] matrix;
	always_comb 
	begin
	R=8'h0;
	G=8'h0;
	B=8'h0;
		pixel = matrix[x][y];
		case(pixel)
		2'd0: begin
			R = 8'h60;
			G = 8'h60;
			B = 8'h60;
		end
		2'd1: begin
			R = 8'd80;
			G = 8'd80;
			B = 8'd80;
		end
		2'd2: begin
			R = 8'd120;
			G = 8'd120;
			B = 8'd120;
		end
		2'd3: begin
			R = 8'd160;
			G = 8'd160;
			B = 8'd160;
		end
		
	endcase
		


matrix = '{
'{2'd0, 2'd0, 2'd0,2'd0,2'd0, 2'd0, 2'd0, 2'd0, 2'd0,2'd0, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2,  2'd2,  2'd2, 2'd2, 2'd2},
'{2'd0, 2'd0, 2'd0,2'd0,2'd0, 2'd0, 2'd0, 2'd0, 2'd0,2'd0, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2,  2'd2,  2'd2, 2'd2, 2'd2},
'{2'd0, 2'd0, 2'd0,2'd0,2'd0, 2'd0, 2'd0, 2'd0, 2'd0,2'd0, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2,  2'd2,  2'd2, 2'd2, 2'd2},
'{2'd0, 2'd0, 2'd0,2'd0,2'd0, 2'd0, 2'd0, 2'd0, 2'd0,2'd0, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2,  2'd2,  2'd2, 2'd2, 2'd2},
'{2'd0, 2'd0, 2'd0,2'd0,2'd0, 2'd0, 2'd0, 2'd0, 2'd0,2'd0, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2,  2'd2,  2'd2, 2'd2, 2'd2},
'{2'd0, 2'd0, 2'd0,2'd0,2'd0, 2'd0, 2'd0, 2'd0, 2'd0,2'd0, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2,  2'd2,  2'd2, 2'd2, 2'd2},
'{2'd0, 2'd0, 2'd0,2'd0,2'd0, 2'd0, 2'd0, 2'd0, 2'd0,2'd0, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2,  2'd2,  2'd2, 2'd2, 2'd2},
'{2'd0, 2'd0, 2'd0,2'd0,2'd0, 2'd0, 2'd0, 2'd0, 2'd0,2'd0, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2,  2'd2,  2'd2, 2'd2, 2'd2},
'{2'd0, 2'd0, 2'd0,2'd0,2'd0, 2'd0, 2'd0, 2'd0, 2'd0,2'd0, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2,  2'd2,  2'd2, 2'd2, 2'd2},
'{2'd0, 2'd0, 2'd0,2'd0,2'd0, 2'd0, 2'd0, 2'd0, 2'd0,2'd0, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2, 2'd2,  2'd2,  2'd2, 2'd2, 2'd2},
'{2'd1, 2'd1, 2'd1,2'd1,2'd1, 2'd1, 2'd1, 2'd1, 2'd1,2'd1, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3,  2'd3,  2'd3, 2'd3, 2'd3},
'{2'd1, 2'd1, 2'd1,2'd1,2'd1, 2'd1, 2'd1, 2'd1, 2'd1,2'd1, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3,  2'd3,  2'd3, 2'd3, 2'd3},
'{2'd1, 2'd1, 2'd1,2'd1,2'd1, 2'd1, 2'd1, 2'd1, 2'd1,2'd1, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3,  2'd3,  2'd3, 2'd3, 2'd3},
'{2'd1, 2'd1, 2'd1,2'd1,2'd1, 2'd1, 2'd1, 2'd1, 2'd1,2'd1, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3,  2'd3,  2'd3, 2'd3, 2'd3},
'{2'd1, 2'd1, 2'd1,2'd1,2'd1, 2'd1, 2'd1, 2'd1, 2'd1,2'd1, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3,  2'd3,  2'd3, 2'd3, 2'd3},
'{2'd1, 2'd1, 2'd1,2'd1,2'd1, 2'd1, 2'd1, 2'd1, 2'd1,2'd1, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3,  2'd3,  2'd3, 2'd3, 2'd3},
'{2'd1, 2'd1, 2'd1,2'd1,2'd1, 2'd1, 2'd1, 2'd1, 2'd1,2'd1, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3,  2'd3,  2'd3, 2'd3, 2'd3},
'{2'd1, 2'd1, 2'd1,2'd1,2'd1, 2'd1, 2'd1, 2'd1, 2'd1,2'd1, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3,  2'd3,  2'd3, 2'd3, 2'd3},
'{2'd1, 2'd1, 2'd1,2'd1,2'd1, 2'd1, 2'd1, 2'd1, 2'd1,2'd1, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3,  2'd3,  2'd3, 2'd3, 2'd3},
'{2'd1, 2'd1, 2'd1,2'd1,2'd1, 2'd1, 2'd1, 2'd1, 2'd1,2'd1, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3, 2'd3,  2'd3,  2'd3, 2'd3, 2'd3}
};
end
endmodule