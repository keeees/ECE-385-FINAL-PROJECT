module background(
					input [9:0] x,
					input [9:0] y,
					output logic [7:0] R,
					output logic [7:0] G,
					output logic [7:0] B
						);
	logic [2:0] pixel;
	//logic [0:][0:499][0:2] matrix;
	logic [0:9][0:9][0:2] matrix;
	always_comb 
	begin
	R=8'h0;
	G=8'h0;
	B=8'h0;
		pixel = matrix[x][y];
		case(pixel)
		3'd0: begin
			R = 8'h0;
			G = 8'h0;
			B = 8'h0;
		end
		3'd1: begin
			R = 8'd11;
			G = 8'd11;
			B = 8'd11;
		end
		3'd2: begin
			R = 8'd100;
			G = 8'd100;
			B = 8'd100;
		end
		3'd3: begin
			R = 8'd120;
			G = 8'd120;
			B = 8'd120;
		end
		3'd4: begin
			R = 8'd90;
			G = 8'd90;
			B = 8'd90;
		end
		3'd5: begin
			R = 8'd95;
			G = 8'd95;
			B = 8'd95;
		end
		3'd6: begin
			R = 8'd105;
			G = 8'd105;
			B = 8'd105;
		end

	endcase
		


matrix = '{
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd0, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd5, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd4, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd0, 3'd6, 3'd1, 3'd0, 3'd1, 3'd5, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0},
'{3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd6, 3'd4, 3'd0, 3'd1, 3'd5, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0}

};
end
endmodule