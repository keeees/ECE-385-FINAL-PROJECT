//
// sawn Wave ROM Table
//
module sawn_table(
  input [7:0] index,
  output [15:0] signal
);
parameter PERIOD = 256; // length of table

assign signal = sawn;
logic [15:0] sawn;
        
always_ff @(index)
begin
case(index)
	8'h00: sawn = 16'h3fff ;
	8'h01: sawn = 16'h3fdf ;
	8'h02: sawn = 16'h3ebf ;
	8'h03: sawn = 16'h3e9f ;
	8'h04: sawn = 16'h3d7f ;
	8'h05: sawn = 16'h3d5f ;
	8'h06: sawn = 16'h3c3f ;
	8'h07: sawn = 16'h3c1f ;
	8'h08: sawn = 16'h3bff ;
	8'h09: sawn = 16'h3bdf ;
	8'h0a: sawn = 16'h3abf ;
	8'h0b: sawn = 16'h3a9f ;
	8'h0c: sawn = 16'h397f ;
	8'h0d: sawn = 16'h395f ;
	8'h0e: sawn = 16'h383f ;
	8'h0f: sawn = 16'h381f ;
	8'h10: sawn = 16'h37ff ;
	8'h11: sawn = 16'h37df ;
	8'h12: sawn = 16'h36bf ;
	8'h13: sawn = 16'h369f ;
	8'h14: sawn = 16'h357f ;
	8'h15: sawn = 16'h355f ;
	8'h16: sawn = 16'h343f ;
	8'h17: sawn = 16'h341f ;
	8'h18: sawn = 16'h33ff ;
	8'h19: sawn = 16'h33df ;
	8'h1a: sawn = 16'h32bf ;
	8'h1b: sawn = 16'h329f ;
	8'h1c: sawn = 16'h317f ;
	8'h1d: sawn = 16'h315f ;
	8'h1e: sawn = 16'h303f ;
	8'h1f: sawn = 16'h301f ;
	8'h20: sawn = 16'h2fff ;
	8'h21: sawn = 16'h2fdf ;
	8'h22: sawn = 16'h2ebf ;
	8'h23: sawn = 16'h2e9f ;
	8'h24: sawn = 16'h2d7f ;
	8'h25: sawn = 16'h2d5f ;
	8'h26: sawn = 16'h2c3f ;
	8'h27: sawn = 16'h2c1f ;
	8'h28: sawn = 16'h2bff ;
	8'h29: sawn = 16'h2bdf ;
	8'h2a: sawn = 16'h2abf ;
	8'h2b: sawn = 16'h2a9f ;
	8'h2c: sawn = 16'h297f ;
	8'h2d: sawn = 16'h295f ;
	8'h2e: sawn = 16'h283f ;
	8'h2f: sawn = 16'h281f ;
	8'h30: sawn = 16'h27ff ;
	8'h31: sawn = 16'h27df ;
	8'h32: sawn = 16'h26bf ;
	8'h33: sawn = 16'h269f ;
	8'h34: sawn = 16'h257f ;
	8'h35: sawn = 16'h255f ;
	8'h36: sawn = 16'h243f ;
	8'h37: sawn = 16'h241f ;
	8'h38: sawn = 16'h23ff ;
	8'h39: sawn = 16'h23df ;
	8'h3a: sawn = 16'h22bf ;
	8'h3b: sawn = 16'h229f ;
	8'h3c: sawn = 16'h217f ;
	8'h3d: sawn = 16'h215f ;
	8'h3e: sawn = 16'h203f ;
	8'h3f: sawn = 16'h201f ;
	8'h40: sawn = 16'h1fff ;
	8'h41: sawn = 16'h1fdf ;
	8'h42: sawn = 16'h1ebf ;
	8'h43: sawn = 16'h1e9f ;
	8'h44: sawn = 16'h1d7f ;
	8'h45: sawn = 16'h1d5f ;
	8'h46: sawn = 16'h1c3f ;
	8'h47: sawn = 16'h1c1f ;
	8'h48: sawn = 16'h1bff ;
	8'h49: sawn = 16'h1bdf ;
	8'h4a: sawn = 16'h1abf ;
	8'h4b: sawn = 16'h1a9f ;
	8'h4c: sawn = 16'h197f ;
	8'h4d: sawn = 16'h195f ;
	8'h4e: sawn = 16'h183f ;
	8'h4f: sawn = 16'h181f ;
	8'h50: sawn = 16'h17ff ;
	8'h51: sawn = 16'h17df ;
	8'h52: sawn = 16'h16bf ;
	8'h53: sawn = 16'h169f ;
	8'h54: sawn = 16'h157f ;
	8'h55: sawn = 16'h155f ;
	8'h56: sawn = 16'h143f ;
	8'h57: sawn = 16'h141f ;
	8'h58: sawn = 16'h13ff ;
	8'h59: sawn = 16'h13df ;
	8'h5a: sawn = 16'h12bf ;
	8'h5b: sawn = 16'h129f ;
	8'h5c: sawn = 16'h117f ;
	8'h5d: sawn = 16'h115f ;
	8'h5e: sawn = 16'h103f ;
	8'h5f: sawn = 16'h101f ;
	8'h60: sawn = 16'h0fff ;
	8'h61: sawn = 16'h0fdf ;
	8'h62: sawn = 16'h0ebf ;
	8'h63: sawn = 16'h0e9f ;
	8'h64: sawn = 16'h0d7f ;
	8'h65: sawn = 16'h0d5f ;
	8'h66: sawn = 16'h0c3f ;
	8'h67: sawn = 16'h0c1f ;
	8'h68: sawn = 16'h0bff ;
	8'h69: sawn = 16'h0bdf ;
	8'h6a: sawn = 16'h0abf ;
	8'h6b: sawn = 16'h0a9f ;
	8'h6c: sawn = 16'h097f ;
	8'h6d: sawn = 16'h095f ;
	8'h6e: sawn = 16'h083f ;
	8'h6f: sawn = 16'h081f ;
	8'h70: sawn = 16'h07ff ;
	8'h71: sawn = 16'h07df ;
	8'h72: sawn = 16'h06bf ;
	8'h73: sawn = 16'h069f ;
	8'h74: sawn = 16'h057f ;
	8'h75: sawn = 16'h0f5f ;
	8'h76: sawn = 16'h053f ;
	8'h77: sawn = 16'h041f ;
	8'h78: sawn = 16'h04ff ;
	8'h79: sawn = 16'h03df ;
	8'h7a: sawn = 16'h03bf ;
	8'h7b: sawn = 16'h029f ;
	8'h7c: sawn = 16'h027f ;
	8'h7d: sawn = 16'h015f ;
	8'h7e: sawn = 16'h013f ;
	8'h7f: sawn = 16'h001f ;
	8'h80: sawn = 16'h0000 ;
	8'h81: sawn = 16'hffe1 ;
	8'h82: sawn = 16'hffc1 ;
	8'h83: sawn = 16'hfea1 ;
	8'h84: sawn = 16'hfe81 ;
	8'h85: sawn = 16'hfd61 ;
	8'h86: sawn = 16'hfd41 ;
	8'h87: sawn = 16'hfc21 ;
	8'h88: sawn = 16'hfc01 ;
	8'h89: sawn = 16'hfbe1 ;
	8'h8a: sawn = 16'hfbc1 ;
	8'h8b: sawn = 16'hfaa1 ;
	8'h8c: sawn = 16'hfa81 ;
	8'h8d: sawn = 16'hf961 ;
	8'h8e: sawn = 16'hf941 ;
	8'h8f: sawn = 16'hf821 ;
	8'h90: sawn = 16'hf801 ;
	8'h91: sawn = 16'hf7e1 ;
	8'h92: sawn = 16'hf7c1 ;
	8'h93: sawn = 16'hf6a1 ;
	8'h94: sawn = 16'hf681 ;
	8'h95: sawn = 16'hf561 ;
	8'h96: sawn = 16'hf541 ;
	8'h97: sawn = 16'hf421 ;
	8'h98: sawn = 16'hf401 ;
	8'h99: sawn = 16'hf3e1 ;
	8'h9a: sawn = 16'hf3c1 ;
	8'h9b: sawn = 16'hf2a1 ;
	8'h9c: sawn = 16'hf281 ;
	8'h9d: sawn = 16'hf161 ;
	8'h9e: sawn = 16'hf141 ;
	8'h9f: sawn = 16'hf021 ;
	8'ha0: sawn = 16'hf001 ;
	8'ha1: sawn = 16'hefe1 ;
	8'ha2: sawn = 16'hefc1 ;
	8'ha3: sawn = 16'heea1 ;
	8'ha4: sawn = 16'hee81 ;
	8'ha5: sawn = 16'hed61 ;
	8'ha6: sawn = 16'hed41 ;
	8'ha7: sawn = 16'hec21 ;
	8'ha8: sawn = 16'hec01 ;
	8'ha9: sawn = 16'hebe1 ;
	8'haa: sawn = 16'hebc1 ;
	8'hab: sawn = 16'heaa1 ;
	8'hac: sawn = 16'hea81 ;
	8'had: sawn = 16'he961 ;
	8'hae: sawn = 16'he941 ;
	8'haf: sawn = 16'he821 ;
	8'hb0: sawn = 16'he801 ;
	8'hb1: sawn = 16'he7e1 ;
	8'hb2: sawn = 16'he7c1 ;
	8'hb3: sawn = 16'he6a1 ;
	8'hb4: sawn = 16'he681 ;
	8'hb5: sawn = 16'he561 ;
	8'hb6: sawn = 16'he541 ;
	8'hb7: sawn = 16'he421 ;
	8'hb8: sawn = 16'he401 ;
	8'hb9: sawn = 16'he3e1 ;
	8'hba: sawn = 16'he3c1 ;
	8'hbb: sawn = 16'he2a1 ;
	8'hbc: sawn = 16'he281 ;
	8'hbd: sawn = 16'he161 ;
	8'hbe: sawn = 16'he141 ;
	8'hbf: sawn = 16'he021 ;
	8'hc0: sawn = 16'he001 ;
	8'hc1: sawn = 16'hdfe1 ;
	8'hc2: sawn = 16'hdfc1 ;
	8'hc3: sawn = 16'hdea1 ;
	8'hc4: sawn = 16'hde81 ;
	8'hc5: sawn = 16'hdd61 ;
	8'hc6: sawn = 16'hdd41 ;
	8'hc7: sawn = 16'hdc21 ;
	8'hc8: sawn = 16'hdc01 ;
	8'hc9: sawn = 16'hdbe1 ;
	8'hca: sawn = 16'hdbc1 ;
	8'hcb: sawn = 16'hdaa1 ;
	8'hcc: sawn = 16'hda81 ;
	8'hcd: sawn = 16'hd961 ;
	8'hce: sawn = 16'hd941 ;
	8'hcf: sawn = 16'hd821 ;
	8'hd0: sawn = 16'hd801 ;
	8'hd1: sawn = 16'hd7e1 ;
	8'hd2: sawn = 16'hd7c1 ;
	8'hd3: sawn = 16'hd6a1 ;
	8'hd4: sawn = 16'hd681 ;
	8'hd5: sawn = 16'hd561 ;
	8'hd6: sawn = 16'hd541 ;
	8'hd7: sawn = 16'hd421 ;
	8'hd8: sawn = 16'hd401 ;
	8'hd9: sawn = 16'hd3e1 ;
	8'hda: sawn = 16'hd3c1 ;
	8'hdb: sawn = 16'hd2a1 ;
	8'hdc: sawn = 16'hd281 ;
	8'hdd: sawn = 16'hd161 ;
	8'hde: sawn = 16'hd141 ;
	8'hdf: sawn = 16'hd021 ;
	8'he0: sawn = 16'hc001 ;
	8'he1: sawn = 16'hcfe1 ;
	8'he2: sawn = 16'hcfc1 ;
	8'he3: sawn = 16'hcea1 ;
	8'he4: sawn = 16'hce81 ;
	8'he5: sawn = 16'hcd61 ;
	8'he6: sawn = 16'hcd41 ;
	8'he7: sawn = 16'hcc21 ;
	8'he8: sawn = 16'hcc01 ;
	8'he9: sawn = 16'hcbe1 ;
	8'hea: sawn = 16'hcbc1 ;
	8'heb: sawn = 16'hcaa1 ;
	8'hec: sawn = 16'hca81 ;
	8'hed: sawn = 16'hc961 ;
	8'hee: sawn = 16'hc941 ;
	8'hef: sawn = 16'hc821 ;
	8'hf0: sawn = 16'hc801 ;
	8'hf1: sawn = 16'hc7e1 ;
	8'hf2: sawn = 16'hc7c1 ;
	8'hf3: sawn = 16'hc6a1 ;
	8'hf4: sawn = 16'hc681 ;
	8'hf5: sawn = 16'hc561 ;
	8'hf6: sawn = 16'hc541 ;
	8'hf7: sawn = 16'hc421 ;
	8'hf8: sawn = 16'hc401 ;
	8'hf9: sawn = 16'hc3e1 ;
	8'hfa: sawn = 16'hc3c1 ;
	8'hfb: sawn = 16'hc2a1 ;
	8'hfc: sawn = 16'hc281 ;
	8'hfd: sawn = 16'hc161 ;
	8'hfe: sawn = 16'hc141 ;
	8'hff: sawn = 16'hc021 ;
	default: sawn = 16'h0000;
endcase
end
endmodule
