//-------------------------------------------------------------------------
//    Color_Mapper.sv                                                    --
//    Stephen Kempf                                                      --
//    3-1-06                                                             --
//                                                                       --
//    Modified by David Kesler  07-16-2008                               --
//    Translated by Joe Meng    07-07-2013                               --
//    Modified by Po-Han Huang  10-06-2017                               --
//                                                                       --
//    Fall 2017 Distribution                                             --
//                                                                       --
//    For use with ECE 385 Lab 8                                         --
//    University of Illinois ECE Department                              --
//-------------------------------------------------------------------------

// color_mapper: Decide which color to be output to VGA for each pixel.
module  color_mapper ( input              is_ball,            // Whether current pixel belongs to ball 
							  input 			is_rball[0:15],				//   or background (computed in ball.sv)
							  //input 			is_rball,
                       input        [9:0] DrawX, DrawY,       // Current pixel coordinates
                       output logic [7:0] VGA_R, VGA_G, VGA_B // VGA RGB output
                     );
    
    logic [7:0] Red, Green, Blue;
    parameter [9:0] Ball_X_Center=320;  // Center position on the X axis

    // Output colors to VGA
    assign VGA_R = Red;
    assign VGA_G = Green;
    assign VGA_B = Blue;
    
    // Assign color based on is_ball signal
    always_comb
    begin
        if (is_ball == 1'b1) 
        begin
            // White ball
            Red = 8'hff;
            Green = 8'hff;
            Blue = 8'hff;
        end
//		  else if(is_rball == 1'b1)
//		  begin
//				Red = 8'hff;
//            Green = 8'h00;
//            Blue = 8'h00;
//		  end
		  else if(is_rball[0] == 1'b1)
		  begin
				Red = 8'h00;
            Green = 8'h00;
            Blue = 8'h00;
		  end
		  else if(is_rball[1] == 1'b1)
		  begin
				Red = 8'h00;
            Green = 8'h00;
            Blue = 8'hff;
		  end
		  else if(is_rball[2] == 1'b1)
		  begin
				Red = 8'h00;
            Green = 8'hff;
            Blue = 8'h00;
		  end

		  else if(is_rball[3] == 1'b1)
		  begin
				Red = 8'h00;
            Green = 8'hff;
            Blue = 8'hff;
		  end
		  else if(is_rball[4] == 1'b1)
		  begin
				Red = 8'hff;
            Green = 8'h00;
            Blue = 8'h00;
		  end
		  else if(is_rball[5] == 1'b1)
		  begin
				Red = 8'hff;
            Green = 8'h00;
            Blue = 8'hff;
		  end
		  else if(is_rball[6] == 1'b1)
		  begin
				Red = 8'hff;
            Green = 8'hff;
            Blue = 8'hff;
		  end
		  else if(is_rball[7] == 1'b1)
		  begin
				Red = 8'hff;
            Green = 8'hff;
            Blue = 8'hff;
		  end
		  else if(is_rball[8] == 1'b1)
		  begin
				Red = 8'h00;
            Green = 8'h00;
            Blue = 8'h00;
		  end
		  else if(is_rball[9] == 1'b1)
		  begin
				Red = 8'h00;
            Green = 8'h00;
            Blue = 8'h00;
		  end
		  else if(is_rball[10] == 1'b1)
		  begin
				Red = 8'h00;
            Green = 8'h00;
            Blue = 8'h00;
		  end
		  else if(is_rball[11] == 1'b1)
		  begin
				Red = 8'h00;
            Green = 8'h00;
            Blue = 8'h00;
		  end
		  else if(is_rball[12] == 1'b1)
		  begin
				Red = 8'h00;
            Green = 8'h00;
            Blue = 8'h00;
		  end
		  else if(is_rball[13] == 1'b1)
		  begin
				Red = 8'h00;
            Green = 8'h00;
            Blue = 8'h00;
		  end
		  else if(is_rball[14] == 1'b1)
		  begin
				Red = 8'h00;
            Green = 8'h00;
            Blue = 8'h00;
		  end
		  else if(is_rball[15] == 1'b1)
		  begin
				Red = 8'h00;
            Green = 8'h00;
            Blue = 8'h00;
		  end
        else 
        begin
            // Background with nice color gradient
            Red = 8'h3f; 
            Green = 8'h00;
            Blue = 8'h7f - {1'b0, DrawX[9:3]};
        end
    end 
    
endmodule
